`timescale 1ns/1ps

module ClkDiv_tb;

/////////////////////////////////////////////////////////
///////////////////// Parameters ////////////////////////
/////////////////////////////////////////////////////////
parameter period = 5;

/////////////////////////////////////////////////////////
///////////////////// Declaratios ///////////////////////
/////////////////////////////////////////////////////////

reg       i_ref_en_tb;
reg       i_rst_n_tb;
reg       i_clk_en_tb;
reg [2:0] i_div_ratio_tb;
wire      o_div_clk_tb;

/////////////////////////////////////////////////////////
///////////////////// Instantiation /////////////////////
/////////////////////////////////////////////////////////

ClkDiv DUT(i_ref_en_tb, i_rst_n_tb, i_clk_en_tb, i_div_ratio_tb, o_div_clk_tb);

/////////////////////////////////////////////////////////
///////////////////// Clock generation //////////////////
/////////////////////////////////////////////////////////

always #(0.5*period) i_ref_en_tb = ~i_ref_en_tb;

/////////////////////////////////////////////////////////
///////////////////// Initial Block /////////////////////
/////////////////////////////////////////////////////////

initial begin

    //System functions.
    $dumpfile("CLK_DIV.vcd") ;       
    $dumpvars; 

    //initialization.
    init;

    //divBy('b000);
    //divBy('b001);
    //divBy('b010);
    //divBy('b011);
    //divBy('b100);
    divBy('b101);
    //divBy('b110);
    //divBy('b111);

    $stop;
end

/////////////////////////////////////////////////////////
///////////////////// Tasks /////////////////////////////
/////////////////////////////////////////////////////////

/////////////// Signals Initialization //////////////////
task init;
begin
    i_ref_en_tb    = 'b0;
    i_rst_n_tb     = 'b1;
    i_clk_en_tb    = 'b0;
    i_div_ratio_tb = 'b0;
    #(10*period);
end
endtask

//////////////////////// Reset /////////////////////////
task reset;
begin
    i_rst_n_tb     = 'b0;
    #period;
    i_rst_n_tb     = 'b1;
    #period;
end
endtask

////////////////// Change the FREQUENCY ////////////////////
task divBy;
input reg [2:0] ratio;
begin
    i_div_ratio_tb = ratio;
    reset;
    i_clk_en_tb    = 'b1;
    #(20*period);
end
endtask

endmodule